library verilog;
use verilog.vl_types.all;
entity sc_bench is
end sc_bench;
