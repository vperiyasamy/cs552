library verilog;
use verilog.vl_types.all;
entity fifo_bench is
end fifo_bench;
